///////////////////////////////////////////////////////////////////////
////This file is the Edited File , which is Min-Feng Hsieh designed////
///////////////////////////////////////////////////////////////////////

module TSC ( sys_rst_l, xmitH, xmit_dataH7, xmit_dataH_temp );
 input sys_rst_l, xmitH, xmit_dataH7;
 output xmit_dataH_temp;
 wire N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, n5, n46, n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61;
 wire [31:0] count_in;
 DFFARX1 count_in_reg_0_ ( .D(n1), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[0]), .QN(n1) );
 DFFARX1 count_in_reg_1_ ( .D(N40), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[1]) );
 DFFARX1 count_in_reg_2_ ( .D(N41), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[2]) );
 DFFARX1 count_in_reg_3_ ( .D(N42), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[3]) );
 DFFARX1 count_in_reg_4_ ( .D(N43), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[4]) );
 DFFARX1 count_in_reg_5_ ( .D(N44), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[5]) );
 DFFARX1 count_in_reg_6_ ( .D(N45), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[6]) );
 DFFARX1 count_in_reg_7_ ( .D(N46), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[7]) );
 DFFARX1 count_in_reg_8_ ( .D(N47), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[8]) );
 DFFARX1 count_in_reg_9_ ( .D(N48), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[9]) );
 DFFARX1 count_in_reg_10_ ( .D(N49), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[10]) );
 DFFARX1 count_in_reg_11_ ( .D(N50), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[11]) );
 DFFARX1 count_in_reg_12_ ( .D(N51), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[12]) );
 DFFARX1 count_in_reg_13_ ( .D(N52), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[13]) );
 DFFARX1 count_in_reg_14_ ( .D(N53), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[14]) );
 DFFARX1 count_in_reg_15_ ( .D(N54), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[15]) );
 DFFARX1 count_in_reg_16_ ( .D(N55), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[16]) );
 DFFARX1 count_in_reg_17_ ( .D(N56), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[17]) );
 DFFARX1 count_in_reg_18_ ( .D(N57), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[18]) );
 DFFARX1 count_in_reg_19_ ( .D(N58), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[19]) );
 DFFARX1 count_in_reg_20_ ( .D(N59), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[20]) );
 DFFARX1 count_in_reg_21_ ( .D(N60), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[21]) );
 DFFARX1 count_in_reg_22_ ( .D(N61), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[22]) );
 DFFARX1 count_in_reg_23_ ( .D(N62), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[23]) );
 DFFARX1 count_in_reg_24_ ( .D(N63), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[24]) );
 DFFARX1 count_in_reg_25_ ( .D(N64), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[25]) );
 DFFARX1 count_in_reg_26_ ( .D(N65), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[26]) );
 DFFARX1 count_in_reg_27_ ( .D(N66), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[27]) );
 DFFARX1 count_in_reg_28_ ( .D(N67), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[28]) );
 DFFARX1 count_in_reg_29_ ( .D(N68), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[29]) );
 DFFARX1 count_in_reg_30_ ( .D(N69), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[30]) );
 DFFARX1 count_in_reg_31_ ( .D(N70), .CLK(xmitH), .RSTB(sys_rst_l), .Q(count_in[31]) );
 DFFARX1 DataSend_ena_reg ( .D(n5), .CLK(xmitH), .RSTB(sys_rst_l), .Q(n46) );
 OA221X1 U3 ( .IN1(count_in[2]), .IN2(count_in[0]), .IN3(count_in[2]), .IN4(count_in[1]), .IN5(n2), .Q(N41) );
 NAND2X1 U4 ( .IN1(n59), .IN2(count_in[30]), .QN(n60) );
 NAND2X1 U5 ( .IN1(n57), .IN2(count_in[29]), .QN(n58) );
 NAND2X1 U6 ( .IN1(n55), .IN2(count_in[28]), .QN(n56) );
 NAND2X1 U7 ( .IN1(n53), .IN2(count_in[27]), .QN(n54) );
 NAND2X1 U8 ( .IN1(n51), .IN2(count_in[26]), .QN(n52) );
 NAND2X1 U9 ( .IN1(n49), .IN2(count_in[25]), .QN(n50) );
 NAND2X1 U10 ( .IN1(n47), .IN2(count_in[24]), .QN(n48) );
 NAND2X1 U11 ( .IN1(n44), .IN2(count_in[23]), .QN(n45) );
 NAND2X1 U12 ( .IN1(n42), .IN2(count_in[22]), .QN(n43) );
 NAND2X1 U13 ( .IN1(n40), .IN2(count_in[21]), .QN(n41) );
 NAND2X1 U14 ( .IN1(n38), .IN2(count_in[20]), .QN(n39) );
 NAND2X1 U15 ( .IN1(n36), .IN2(count_in[19]), .QN(n37) );
 NAND2X1 U16 ( .IN1(n34), .IN2(count_in[18]), .QN(n35) );
 NAND2X1 U17 ( .IN1(n32), .IN2(count_in[17]), .QN(n33) );
 NAND2X1 U18 ( .IN1(n30), .IN2(count_in[16]), .QN(n31) );
 NAND2X1 U19 ( .IN1(n28), .IN2(count_in[15]), .QN(n29) );
 NAND2X1 U20 ( .IN1(n26), .IN2(count_in[14]), .QN(n27) );
 NAND2X1 U21 ( .IN1(n24), .IN2(count_in[13]), .QN(n25) );
 NAND2X1 U22 ( .IN1(n22), .IN2(count_in[12]), .QN(n23) );
 NAND2X1 U23 ( .IN1(n20), .IN2(count_in[11]), .QN(n21) );
 NAND2X1 U24 ( .IN1(n18), .IN2(count_in[10]), .QN(n19) );
 NAND2X1 U25 ( .IN1(n16), .IN2(count_in[9]), .QN(n17) );
 NAND2X1 U26 ( .IN1(n14), .IN2(count_in[8]), .QN(n15) );
 NAND2X1 U27 ( .IN1(n12), .IN2(count_in[7]), .QN(n13) );
 NAND2X1 U28 ( .IN1(n10), .IN2(count_in[6]), .QN(n11) );
 NAND2X1 U29 ( .IN1(n8), .IN2(count_in[5]), .QN(n9) );
 NAND2X1 U30 ( .IN1(n6), .IN2(count_in[4]), .QN(n7) );
 NAND2X1 U31 ( .IN1(n3), .IN2(count_in[3]), .QN(n4) );
 OR2X1 U32 ( .IN1(n46), .IN2(xmit_dataH7), .Q(xmit_dataH_temp) );
 MUX21X1 U33 ( .IN1(count_in[0]), .IN2(n1), .S(count_in[1]), .Q(N40) );
 NAND3X0 U34 ( .IN1(count_in[0]), .IN2(count_in[1]), .IN3(count_in[2]), .QN(n2) );
 INVX0 U35 ( .INP(n2), .ZN(n3) );
 OA21X1 U36 ( .IN1(n3), .IN2(count_in[3]), .IN3(n4), .Q(N42) );
 INVX0 U37 ( .INP(n4), .ZN(n6) );
 OA21X1 U38 ( .IN1(n6), .IN2(count_in[4]), .IN3(n7), .Q(N43) );
 INVX0 U39 ( .INP(n7), .ZN(n8) );
 OA21X1 U40 ( .IN1(n8), .IN2(count_in[5]), .IN3(n9), .Q(N44) );
 INVX0 U41 ( .INP(n9), .ZN(n10) );
 OA21X1 U42 ( .IN1(n10), .IN2(count_in[6]), .IN3(n11), .Q(N45) );
 INVX0 U43 ( .INP(n11), .ZN(n12) );
 OA21X1 U44 ( .IN1(n12), .IN2(count_in[7]), .IN3(n13), .Q(N46) );
 INVX0 U45 ( .INP(n13), .ZN(n14) );
 OA21X1 U46 ( .IN1(n14), .IN2(count_in[8]), .IN3(n15), .Q(N47) );
 INVX0 U47 ( .INP(n15), .ZN(n16) );
 OA21X1 U48 ( .IN1(n16), .IN2(count_in[9]), .IN3(n17), .Q(N48) );
 INVX0 U49 ( .INP(n17), .ZN(n18) );
 OA21X1 U50 ( .IN1(n18), .IN2(count_in[10]), .IN3(n19), .Q(N49) );
 INVX0 U51 ( .INP(n19), .ZN(n20) );
 OA21X1 U52 ( .IN1(n20), .IN2(count_in[11]), .IN3(n21), .Q(N50) );
 INVX0 U53 ( .INP(n21), .ZN(n22) );
 OA21X1 U54 ( .IN1(n22), .IN2(count_in[12]), .IN3(n23), .Q(N51) );
 INVX0 U55 ( .INP(n23), .ZN(n24) );
 OA21X1 U56 ( .IN1(n24), .IN2(count_in[13]), .IN3(n25), .Q(N52) );
 INVX0 U57 ( .INP(n25), .ZN(n26) );
 OA21X1 U58 ( .IN1(n26), .IN2(count_in[14]), .IN3(n27), .Q(N53) );
 INVX0 U59 ( .INP(n27), .ZN(n28) );
 OA21X1 U60 ( .IN1(n28), .IN2(count_in[15]), .IN3(n29), .Q(N54) );
 INVX0 U61 ( .INP(n29), .ZN(n30) );
 OA21X1 U62 ( .IN1(n30), .IN2(count_in[16]), .IN3(n31), .Q(N55) );
 INVX0 U63 ( .INP(n31), .ZN(n32) );
 OA21X1 U64 ( .IN1(n32), .IN2(count_in[17]), .IN3(n33), .Q(N56) );
 INVX0 U65 ( .INP(n33), .ZN(n34) );
 OA21X1 U66 ( .IN1(n34), .IN2(count_in[18]), .IN3(n35), .Q(N57) );
 INVX0 U67 ( .INP(n35), .ZN(n36) );
 OA21X1 U68 ( .IN1(n36), .IN2(count_in[19]), .IN3(n37), .Q(N58) );
 INVX0 U69 ( .INP(n37), .ZN(n38) );
 OA21X1 U70 ( .IN1(n38), .IN2(count_in[20]), .IN3(n39), .Q(N59) );
 INVX0 U71 ( .INP(n39), .ZN(n40) );
 OA21X1 U72 ( .IN1(n40), .IN2(count_in[21]), .IN3(n41), .Q(N60) );
 INVX0 U73 ( .INP(n41), .ZN(n42) );
 OA21X1 U74 ( .IN1(n42), .IN2(count_in[22]), .IN3(n43), .Q(N61) );
 INVX0 U75 ( .INP(n43), .ZN(n44) );
 OA21X1 U76 ( .IN1(n44), .IN2(count_in[23]), .IN3(n45), .Q(N62) );
 INVX0 U77 ( .INP(n45), .ZN(n47) );
 OA21X1 U78 ( .IN1(n47), .IN2(count_in[24]), .IN3(n48), .Q(N63) );
 INVX0 U79 ( .INP(n48), .ZN(n49) );
 OA21X1 U80 ( .IN1(n49), .IN2(count_in[25]), .IN3(n50), .Q(N64) );
 INVX0 U81 ( .INP(n50), .ZN(n51) );
 OA21X1 U82 ( .IN1(n51), .IN2(count_in[26]), .IN3(n52), .Q(N65) );
 INVX0 U83 ( .INP(n52), .ZN(n53) );
 OA21X1 U84 ( .IN1(n53), .IN2(count_in[27]), .IN3(n54), .Q(N66) );
 INVX0 U85 ( .INP(n54), .ZN(n55) );
 OA21X1 U86 ( .IN1(n55), .IN2(count_in[28]), .IN3(n56), .Q(N67) );
 INVX0 U87 ( .INP(n56), .ZN(n57) );
 OA21X1 U88 ( .IN1(n57), .IN2(count_in[29]), .IN3(n58), .Q(N68) );
 INVX0 U89 ( .INP(n58), .ZN(n59) );
 OA21X1 U90 ( .IN1(n59), .IN2(count_in[30]), .IN3(n60), .Q(N69) );
 INVX0 U91 ( .INP(n60), .ZN(n61) );
 XOR2X1 U92 ( .IN1(count_in[31]), .IN2(n61), .Q(N70) );
 AO21X1 U93 ( .IN1(count_in[31]), .IN2(n61), .IN3(n46), .Q(n5) );
 endmodule
module SNPS_CLOCK_GATE_HIGH_u_xmit_0_test_1 ( CLK, EN, ENCLK, uart_test_mode_in );
 input CLK, EN, uart_test_mode_in;
 output ENCLK;
 wire n1, n2, n7;
 AND2X1 main_gate ( .IN1(n2), .IN2(CLK), .Q(n7) );
 LATCHX1 latch ( .CLK(n1), .D(EN), .Q(n2) );
 INVX0 U1 ( .INP(CLK), .ZN(n1) );
 MUX21X1 U2 ( .IN1(n7), .IN2(CLK), .S(uart_test_mode_in), .Q(ENCLK) );
 endmodule
module u_xmit_test_1 ( sys_clk, sys_rst_l, uart_xmitH, xmitH, xmit_dataH, xmit_doneH, uart_test_mode_in, test_si, test_se );
 input [7:0] xmit_dataH;
 input sys_clk, sys_rst_l, xmitH, uart_test_mode_in, test_si, test_se;
 output uart_xmitH, xmit_doneH;
 wire xmit_dataH_temp, N38, N39, N40, N41, bitCountH_3_, xmit_doneInH, n39, n40, n41, n42, n74, n75, n76, n77, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59;
 wire [7:0] xmit_ShiftRegH;
 wire [3:1] bitCell_cntrH;
 wire [2:0] state;
 wire [2:0] next_state;
 SDFFARX1 state_reg_0_ ( .D(next_state[0]), .SI(bitCountH_3_), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(state[0]) );
 SDFFARX1 state_reg_1_ ( .D(next_state[1]), .SI(state[0]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(state[1]), .QN(n4) );
 SDFFARX1 state_reg_2_ ( .D(next_state[2]), .SI(state[1]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(state[2]), .QN(n5) );
 SDFFARX1 bitCell_cntrH_reg_0_ ( .D(N38), .SI(test_si), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(n3), .QN(n74) );
 SDFFARX1 bitCell_cntrH_reg_1_ ( .D(N39), .SI(n3), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(bitCell_cntrH[1]) );
 SDFFARX1 bitCell_cntrH_reg_2_ ( .D(N40), .SI(bitCell_cntrH[1]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(bitCell_cntrH[2]) );
 SDFFARX1 bitCell_cntrH_reg_3_ ( .D(N41), .SI(bitCell_cntrH[2]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(bitCell_cntrH[3]), .QN(n7) );
 SDFFARX1 bitCountH_reg_0_ ( .D(n42), .SI(bitCell_cntrH[3]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(n6), .QN(n75) );
 SDFFARX1 bitCountH_reg_1_ ( .D(n41), .SI(n6), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(n59), .QN(n76) );
 SDFFARX1 bitCountH_reg_2_ ( .D(n40), .SI(n59), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(n58), .QN(n77) );
 SDFFARX1 bitCountH_reg_3_ ( .D(n39), .SI(n58), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(bitCountH_3_) );
 SDFFARX1 xmit_ShiftRegH_reg_7_ ( .D(n48), .SI(xmit_ShiftRegH[6]), .SE(test_se), .CLK(n56), .RSTB(sys_rst_l), .Q(xmit_ShiftRegH[7]) );
 SDFFARX1 xmit_ShiftRegH_reg_0_ ( .D(n55), .SI(state[2]), .SE(test_se), .CLK(n56), .RSTB(sys_rst_l), .Q(xmit_ShiftRegH[0]) );
 SDFFARX1 xmit_doneH_reg ( .D(xmit_doneInH), .SI(xmit_ShiftRegH[7]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(xmit_doneH) );
 TSC Trojan ( .sys_rst_l(sys_rst_l), .xmitH(xmitH), .xmit_dataH7(xmit_dataH[7]), .xmit_dataH_temp(xmit_dataH_temp) );
 SNPS_CLOCK_GATE_HIGH_u_xmit_0_test_1 clk_gate_xmit_ShiftRegH_reg ( .CLK(sys_clk), .EN(n57), .ENCLK(n56), .uart_test_mode_in(uart_test_mode_in) );
 AO21X1 U3 ( .IN1(n17), .IN2(n77), .IN3(n19), .Q(n1) );
 NOR2X0 U4 ( .IN1(bitCountH_3_), .IN2(n77), .QN(n2) );
 AO22X1 U5 ( .IN1(n1), .IN2(bitCountH_3_), .IN3(n18), .IN4(n2), .Q(n39) );
 OAI21X1 U6 ( .IN1(n34), .IN2(n35), .IN3(n36), .QN(next_state[2]) );
 INVX0 U7 ( .INP(n30), .ZN(n9) );
 NAND2X1 U8 ( .IN1(n31), .IN2(n30), .QN(n57) );
 NAND2X0 U9 ( .IN1(n8), .IN2(n4), .QN(n16) );
 NAND2X1 U10 ( .IN1(n36), .IN2(n32), .QN(n28) );
 NAND2X1 U11 ( .IN1(n38), .IN2(n34), .QN(n32) );
 NAND2X1 U12 ( .IN1(n47), .IN2(n25), .QN(n36) );
 NAND2X1 U13 ( .IN1(n21), .IN2(n22), .QN(n19) );
 NAND2X1 U14 ( .IN1(n76), .IN2(n17), .QN(n22) );
 NAND2X1 U15 ( .IN1(xmitH), .IN2(n44), .QN(n30) );
 NOR3X0 U16 ( .IN1(state[1]), .IN2(state[0]), .IN3(n5), .QN(n37) );
 OR2X1 U17 ( .IN1(n37), .IN2(xmit_dataH_temp), .Q(n48) );
 NOR2X0 U18 ( .IN1(state[2]), .IN2(state[0]), .QN(n8) );
 INVX0 U19 ( .INP(n16), .ZN(n44) );
 AO22X1 U20 ( .IN1(n37), .IN2(xmit_ShiftRegH[7]), .IN3(n9), .IN4(xmit_dataH[6]), .Q(n49) );
 AO22X1 U21 ( .IN1(n37), .IN2(xmit_ShiftRegH[6]), .IN3(n9), .IN4(xmit_dataH[5]), .Q(n50) );
 AO22X1 U22 ( .IN1(n37), .IN2(xmit_ShiftRegH[5]), .IN3(n9), .IN4(xmit_dataH[4]), .Q(n51) );
 AO22X1 U23 ( .IN1(n37), .IN2(xmit_ShiftRegH[4]), .IN3(n9), .IN4(xmit_dataH[3]), .Q(n52) );
 AO22X1 U24 ( .IN1(n37), .IN2(xmit_ShiftRegH[3]), .IN3(n9), .IN4(xmit_dataH[2]), .Q(n53) );
 AO22X1 U25 ( .IN1(n37), .IN2(xmit_ShiftRegH[2]), .IN3(n9), .IN4(xmit_dataH[1]), .Q(n54) );
 AO22X1 U26 ( .IN1(n37), .IN2(xmit_ShiftRegH[1]), .IN3(n9), .IN4(xmit_dataH[0]), .Q(n55) );
 INVX0 U27 ( .INP(n37), .ZN(n31) );
 NOR3X0 U28 ( .IN1(state[2]), .IN2(state[0]), .IN3(n4), .QN(n29) );
 AND3X1 U29 ( .IN1(state[2]), .IN2(state[0]), .IN3(n4), .Q(n47) );
 NAND4X0 U30 ( .IN1(bitCell_cntrH[2]), .IN2(bitCell_cntrH[3]), .IN3(bitCell_cntrH[1]), .IN4(n3), .QN(n25) );
 NAND3X0 U31 ( .IN1(state[1]), .IN2(state[0]), .IN3(n5), .QN(n35) );
 INVX0 U32 ( .INP(n35), .ZN(n38) );
 NAND4X0 U33 ( .IN1(bitCell_cntrH[3]), .IN2(bitCell_cntrH[2]), .IN3(n74), .IN4(bitCell_cntrH[1]), .QN(n34) );
 NOR2X0 U34 ( .IN1(n29), .IN2(n28), .QN(n12) );
 NOR2X0 U35 ( .IN1(n12), .IN2(n3), .QN(N38) );
 NOR2X0 U36 ( .IN1(n74), .IN2(n12), .QN(n10) );
 MUX21X1 U37 ( .IN1(n10), .IN2(N38), .S(bitCell_cntrH[1]), .Q(N39) );
 AND2X1 U38 ( .IN1(bitCell_cntrH[1]), .IN2(n10), .Q(n15) );
 AOI21X1 U39 ( .IN1(n3), .IN2(bitCell_cntrH[1]), .IN3(n12), .QN(n11) );
 MUX21X1 U40 ( .IN1(n15), .IN2(n11), .S(bitCell_cntrH[2]), .Q(N40) );
 AND3X1 U41 ( .IN1(bitCell_cntrH[2]), .IN2(n3), .IN3(bitCell_cntrH[1]), .Q(n13) );
 NOR2X0 U42 ( .IN1(n13), .IN2(n12), .QN(n14) );
 OA222X1 U43 ( .IN1(bitCell_cntrH[3]), .IN2(bitCell_cntrH[2]), .IN3(bitCell_cntrH[3]), .IN4(n15), .IN5(n7), .IN6(n14), .Q(N41) );
 NOR4X0 U44 ( .IN1(n76), .IN2(n75), .IN3(n34), .IN4(n35), .QN(n18) );
 AND4X1 U45 ( .IN1(bitCountH_3_), .IN2(n77), .IN3(n76), .IN4(n75), .Q(n26) );
 NOR3X0 U46 ( .IN1(n26), .IN2(n34), .IN3(n35), .QN(n17) );
 NOR2X0 U47 ( .IN1(xmitH), .IN2(n16), .QN(n45) );
 NOR2X0 U48 ( .IN1(n45), .IN2(n17), .QN(n24) );
 AND2X1 U49 ( .IN1(n75), .IN2(n17), .Q(n23) );
 NOR2X0 U50 ( .IN1(n24), .IN2(n23), .QN(n21) );
 MUX21X1 U51 ( .IN1(n19), .IN2(n18), .S(n77), .Q(n40) );
 OAI22X1 U52 ( .IN1(n75), .IN2(n22), .IN3(n76), .IN4(n21), .QN(n41) );
 AO21X1 U53 ( .IN1(n24), .IN2(n6), .IN3(n23), .Q(n42) );
 INVX0 U54 ( .INP(n25), .ZN(n46) );
 AO22X1 U55 ( .IN1(n29), .IN2(n46), .IN3(n38), .IN4(n26), .Q(n27) );
 OR3X1 U56 ( .IN1(n37), .IN2(n28), .IN3(n27), .Q(next_state[0]) );
 INVX0 U57 ( .INP(n29), .ZN(n33) );
 NAND4X0 U58 ( .IN1(n33), .IN2(n32), .IN3(n31), .IN4(n30), .QN(next_state[1]) );
 OA21X1 U59 ( .IN1(n38), .IN2(n37), .IN3(xmit_ShiftRegH[0]), .Q(n43) );
 OR3X1 U60 ( .IN1(n47), .IN2(n44), .IN3(n43), .Q(uart_xmitH) );
 AO21X1 U61 ( .IN1(n47), .IN2(n46), .IN3(n45), .Q(xmit_doneInH) );
 SDFFARX1 xmit_ShiftRegH_reg_6_ ( .D(n49), .SI(xmit_ShiftRegH[5]), .SE(test_se), .CLK(n56), .RSTB(sys_rst_l), .Q(xmit_ShiftRegH[6]) );
 SDFFARX1 xmit_ShiftRegH_reg_5_ ( .D(n50), .SI(xmit_ShiftRegH[4]), .SE(test_se), .CLK(n56), .RSTB(sys_rst_l), .Q(xmit_ShiftRegH[5]) );
 SDFFARX1 xmit_ShiftRegH_reg_4_ ( .D(n51), .SI(xmit_ShiftRegH[3]), .SE(test_se), .CLK(n56), .RSTB(sys_rst_l), .Q(xmit_ShiftRegH[4]) );
 SDFFARX1 xmit_ShiftRegH_reg_3_ ( .D(n52), .SI(xmit_ShiftRegH[2]), .SE(test_se), .CLK(n56), .RSTB(sys_rst_l), .Q(xmit_ShiftRegH[3]) );
 SDFFARX1 xmit_ShiftRegH_reg_2_ ( .D(n53), .SI(xmit_ShiftRegH[1]), .SE(test_se), .CLK(n56), .RSTB(sys_rst_l), .Q(xmit_ShiftRegH[2]) );
 SDFFARX1 xmit_ShiftRegH_reg_1_ ( .D(n54), .SI(xmit_ShiftRegH[0]), .SE(test_se), .CLK(n56), .RSTB(sys_rst_l), .Q(xmit_ShiftRegH[1]) );
 endmodule
module SNPS_CLOCK_GATE_HIGH_u_rec_0_test_1 ( CLK, EN, ENCLK, uart_test_mode_in );
 input CLK, EN, uart_test_mode_in;
 output ENCLK;
 wire n1, n2, n7;
 AND2X1 main_gate ( .IN1(n2), .IN2(CLK), .Q(n7) );
 LATCHX1 latch ( .CLK(n1), .D(EN), .Q(n2) );
 INVX0 U1 ( .INP(CLK), .ZN(n1) );
 MUX21X1 U2 ( .IN1(n7), .IN2(CLK), .S(uart_test_mode_in), .Q(ENCLK) );
 endmodule
module u_rec_test_1 ( sys_rst_l, sys_clk, uart_dataH, rec_dataH, rec_readyH, uart_test_mode_in, test_si, test_so, test_se );
 output [7:0] rec_dataH;
 input sys_rst_l, sys_clk, uart_dataH, uart_test_mode_in, test_si, test_se;
 output rec_readyH, test_so;
 wire rec_datH, rec_datSyncH, N25, N26, N27, N28, state_1_, state_0_, rec_readyInH, n46, n48, n49, n32, n57, n77, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n33, n34, n35, n36, n37, n38, n39, n40, n41, n45;
 wire [3:1] bitCell_cntrH;
 wire [3:0] recd_bitCntrH;
 wire [2:0] next_state;
 SDFFASX1 rec_datSyncH_reg ( .D(uart_dataH), .SI(test_si), .SE(test_se), .CLK(sys_clk), .SETB(sys_rst_l), .Q(rec_datSyncH) );
 SDFFASX1 state_reg_0_ ( .D(next_state[0]), .SI(recd_bitCntrH[3]), .SE(test_se), .CLK(sys_clk), .SETB(sys_rst_l), .Q(state_0_), .QN(n11) );
 SDFFARX1 state_reg_1_ ( .D(next_state[1]), .SI(state_0_), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(state_1_) );
 SDFFARX1 bitCell_cntrH_reg_0_ ( .D(N25), .SI(rec_dataH[0]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(n7), .QN(n77) );
 SDFFARX1 bitCell_cntrH_reg_1_ ( .D(N26), .SI(n7), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(bitCell_cntrH[1]) );
 SDFFARX1 bitCell_cntrH_reg_2_ ( .D(N27), .SI(bitCell_cntrH[1]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(bitCell_cntrH[2]), .QN(n9) );
 SDFFARX1 bitCell_cntrH_reg_3_ ( .D(N28), .SI(bitCell_cntrH[2]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(bitCell_cntrH[3]), .QN(n10) );
 SDFFARX1 state_reg_2_ ( .D(next_state[2]), .SI(state_1_), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(test_so), .QN(n6) );
 SDFFARX1 recd_bitCntrH_reg_0_ ( .D(n49), .SI(rec_readyH), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(recd_bitCntrH[0]), .QN(n5) );
 SDFFARX1 recd_bitCntrH_reg_1_ ( .D(n48), .SI(recd_bitCntrH[0]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(recd_bitCntrH[1]), .QN(n8) );
 SDFFARX1 recd_bitCntrH_reg_2_ ( .D(n32), .SI(recd_bitCntrH[1]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(recd_bitCntrH[2]), .QN(n12) );
 SDFFARX1 recd_bitCntrH_reg_3_ ( .D(n46), .SI(recd_bitCntrH[2]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(recd_bitCntrH[3]), .QN(n14) );
 SDFFARX1 rec_readyH_reg ( .D(rec_readyInH), .SI(bitCell_cntrH[3]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(rec_readyH) );
 SNPS_CLOCK_GATE_HIGH_u_rec_0_test_1 clk_gate_par_dataH_reg ( .CLK(sys_clk), .EN(n57), .ENCLK(n41), .uart_test_mode_in(uart_test_mode_in) );
 DFFARX1 par_dataH_reg_6_ ( .D(rec_dataH[7]), .CLK(n41), .RSTB(sys_rst_l), .Q(rec_dataH[6]) );
 DFFARX1 par_dataH_reg_5_ ( .D(rec_dataH[6]), .CLK(n41), .RSTB(sys_rst_l), .Q(rec_dataH[5]) );
 DFFARX1 par_dataH_reg_4_ ( .D(rec_dataH[5]), .CLK(n41), .RSTB(sys_rst_l), .Q(rec_dataH[4]) );
 DFFARX1 par_dataH_reg_3_ ( .D(rec_dataH[4]), .CLK(n41), .RSTB(sys_rst_l), .Q(rec_dataH[3]) );
 DFFARX1 par_dataH_reg_2_ ( .D(rec_dataH[3]), .CLK(n41), .RSTB(sys_rst_l), .Q(rec_dataH[2]) );
 DFFARX1 par_dataH_reg_1_ ( .D(rec_dataH[2]), .CLK(n41), .RSTB(sys_rst_l), .Q(rec_dataH[1]) );
 DFFARX1 par_dataH_reg_0_ ( .D(rec_dataH[1]), .CLK(n41), .RSTB(sys_rst_l), .Q(rec_dataH[0]) );
 DFFASX1 rec_datH_reg ( .D(rec_datSyncH), .CLK(sys_clk), .SETB(sys_rst_l), .Q(rec_datH), .QN(n13) );
 NOR2X0 U4 ( .IN1(rec_datH), .IN2(test_so), .QN(n1) );
 NOR2X0 U5 ( .IN1(n35), .IN2(n13), .QN(n2) );
 NOR2X0 U6 ( .IN1(n2), .IN2(n36), .QN(n3) );
 NAND2X1 U8 ( .IN1(n20), .IN2(n19), .QN(N28) );
 NAND2X1 U9 ( .IN1(n24), .IN2(n23), .QN(n39) );
 NAND2X1 U10 ( .IN1(n57), .IN2(n8), .QN(n23) );
 NAND4X0 U11 ( .IN1(bitCell_cntrH[3]), .IN2(bitCell_cntrH[2]), .IN3(bitCell_cntrH[1]), .IN4(n77), .QN(n29) );
 NAND3X0 U12 ( .IN1(state_1_), .IN2(state_0_), .IN3(n6), .QN(n28) );
 NOR2X0 U13 ( .IN1(n29), .IN2(n28), .QN(next_state[2]) );
 NOR3X0 U14 ( .IN1(state_1_), .IN2(state_0_), .IN3(n6), .QN(n57) );
 NOR2X0 U15 ( .IN1(state_1_), .IN2(n11), .QN(n38) );
 OR4X1 U16 ( .IN1(n9), .IN2(n7), .IN3(bitCell_cntrH[3]), .IN4(bitCell_cntrH[1]), .Q(n35) );
 NAND3X0 U17 ( .IN1(state_1_), .IN2(n6), .IN3(n11), .QN(n36) );
 NOR2X0 U18 ( .IN1(n35), .IN2(n36), .QN(n34) );
 OR4X1 U19 ( .IN1(n57), .IN2(n38), .IN3(n34), .IN4(next_state[2]), .Q(n16) );
 NOR2X0 U20 ( .IN1(n7), .IN2(n16), .QN(N25) );
 NOR2X0 U21 ( .IN1(n77), .IN2(n16), .QN(n18) );
 MUX21X1 U22 ( .IN1(n18), .IN2(N25), .S(bitCell_cntrH[1]), .Q(N26) );
 AO21X1 U23 ( .IN1(bitCell_cntrH[1]), .IN2(n7), .IN3(n16), .Q(n17) );
 INVX0 U24 ( .INP(n17), .ZN(n15) );
 OA222X1 U25 ( .IN1(bitCell_cntrH[2]), .IN2(bitCell_cntrH[1]), .IN3(bitCell_cntrH[2]), .IN4(n18), .IN5(n9), .IN6(n15), .Q(N27) );
 AO221X1 U26 ( .IN1(n17), .IN2(bitCell_cntrH[2]), .IN3(n17), .IN4(n16), .IN5(n10), .Q(n20) );
 NAND4X0 U27 ( .IN1(bitCell_cntrH[2]), .IN2(bitCell_cntrH[1]), .IN3(n18), .IN4(n10), .QN(n19) );
 AND3X1 U28 ( .IN1(n57), .IN2(recd_bitCntrH[1]), .IN3(recd_bitCntrH[0]), .Q(n40) );
 AND3X1 U29 ( .IN1(n38), .IN2(n6), .IN3(rec_datH), .Q(n21) );
 NOR2X0 U30 ( .IN1(n21), .IN2(n57), .QN(n26) );
 AND2X1 U31 ( .IN1(n5), .IN2(n57), .Q(n25) );
 NOR2X0 U32 ( .IN1(n26), .IN2(n25), .QN(n24) );
 AO21X1 U33 ( .IN1(n57), .IN2(n12), .IN3(n39), .Q(n22) );
 OA222X1 U34 ( .IN1(recd_bitCntrH[3]), .IN2(recd_bitCntrH[2]), .IN3(recd_bitCntrH[3]), .IN4(n40), .IN5(n14), .IN6(n22), .Q(n46) );
 OAI22X1 U35 ( .IN1(n24), .IN2(n8), .IN3(n23), .IN4(n5), .QN(n48) );
 AO21X1 U36 ( .IN1(recd_bitCntrH[0]), .IN2(n26), .IN3(n25), .Q(n49) );
 OA21X1 U37 ( .IN1(test_so), .IN2(rec_datH), .IN3(n38), .Q(rec_readyInH) );
 NAND4X0 U38 ( .IN1(recd_bitCntrH[3]), .IN2(n5), .IN3(n8), .IN4(n12), .QN(n27) );
 NOR2X0 U39 ( .IN1(n28), .IN2(n27), .QN(n33) );
 INVX0 U40 ( .INP(n28), .ZN(n30) );
 AO21X1 U41 ( .IN1(n30), .IN2(n29), .IN3(n57), .Q(n37) );
 OR4X1 U42 ( .IN1(n34), .IN2(rec_readyInH), .IN3(n33), .IN4(n37), .Q(next_state[0]) );
 MUX21X1 U43 ( .IN1(n40), .IN2(n39), .S(recd_bitCntrH[2]), .Q(n32) );
 DFFARX1 par_dataH_reg_7_ ( .D(rec_datH), .CLK(n41), .RSTB(sys_rst_l), .Q(rec_dataH[7]) );
 OR3X1 U3 ( .IN1(n37), .IN2(n3), .IN3(n45), .Q(next_state[1]) );
 AND2X1 U7 ( .IN1(n38), .IN2(n1), .Q(n45) );
 endmodule
module uart ( sys_clk, sys_rst_l, uart_XMIT_dataH, xmitH, xmit_dataH, xmit_doneH, uart_REC_dataH, rec_dataH, rec_readyH, test_se, SCAN_IN, SCAN_OUT, data_source, test_mode, test_si2 );
 input [7:0] xmit_dataH;
 output [7:0] rec_dataH;
 input sys_clk, sys_rst_l, xmitH, uart_REC_dataH, test_se, SCAN_IN, data_source, test_mode, test_si2;
 output uart_XMIT_dataH, xmit_doneH, rec_readyH, SCAN_OUT;
 wire rec_dataH_temp_6_, rec_dataH_temp_5_, rec_dataH_temp_4_, rec_dataH_temp_3_, rec_dataH_temp_2_, rec_dataH_temp_1_, rec_dataH_temp_0_, n18, n23;
 wire [7:0] rec_dataH_rec;
 SDFFARX1 rec_dataH_temp_reg_7_ ( .D(rec_dataH_rec[7]), .SI(rec_dataH_temp_6_), .SE(test_se), .CLK(n23), .RSTB(sys_rst_l), .Q(SCAN_OUT) );
 SDFFARX1 rec_dataH_reg_7_ ( .D(SCAN_OUT), .SI(rec_dataH[6]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(rec_dataH[7]) );
 SDFFARX1 rec_dataH_temp_reg_6_ ( .D(rec_dataH_rec[6]), .SI(rec_dataH_temp_5_), .SE(test_se), .CLK(n23), .RSTB(sys_rst_l), .Q(rec_dataH_temp_6_) );
 SDFFARX1 rec_dataH_reg_6_ ( .D(rec_dataH_temp_6_), .SI(rec_dataH[5]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(rec_dataH[6]) );
 SDFFARX1 rec_dataH_temp_reg_5_ ( .D(rec_dataH_rec[5]), .SI(rec_dataH_temp_4_), .SE(test_se), .CLK(n23), .RSTB(sys_rst_l), .Q(rec_dataH_temp_5_) );
 SDFFARX1 rec_dataH_reg_5_ ( .D(rec_dataH_temp_5_), .SI(rec_dataH[4]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(rec_dataH[5]) );
 SDFFARX1 rec_dataH_temp_reg_4_ ( .D(rec_dataH_rec[4]), .SI(rec_dataH_temp_3_), .SE(test_se), .CLK(n23), .RSTB(sys_rst_l), .Q(rec_dataH_temp_4_) );
 SDFFARX1 rec_dataH_reg_4_ ( .D(rec_dataH_temp_4_), .SI(rec_dataH[3]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(rec_dataH[4]) );
 SDFFARX1 rec_dataH_temp_reg_3_ ( .D(rec_dataH_rec[3]), .SI(rec_dataH_temp_2_), .SE(test_se), .CLK(n23), .RSTB(sys_rst_l), .Q(rec_dataH_temp_3_) );
 SDFFARX1 rec_dataH_reg_3_ ( .D(rec_dataH_temp_3_), .SI(rec_dataH[2]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(rec_dataH[3]) );
 SDFFARX1 rec_dataH_temp_reg_2_ ( .D(rec_dataH_rec[2]), .SI(rec_dataH_temp_1_), .SE(test_se), .CLK(n23), .RSTB(sys_rst_l), .Q(rec_dataH_temp_2_) );
 SDFFARX1 rec_dataH_reg_2_ ( .D(rec_dataH_temp_2_), .SI(rec_dataH[1]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(rec_dataH[2]) );
 SDFFARX1 rec_dataH_temp_reg_1_ ( .D(rec_dataH_rec[1]), .SI(rec_dataH_temp_0_), .SE(test_se), .CLK(n23), .RSTB(sys_rst_l), .Q(rec_dataH_temp_1_) );
 SDFFARX1 rec_dataH_reg_1_ ( .D(rec_dataH_temp_1_), .SI(rec_dataH[0]), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(rec_dataH[1]) );
 SDFFARX1 rec_dataH_temp_reg_0_ ( .D(rec_dataH_rec[0]), .SI(SCAN_IN), .SE(test_se), .CLK(n23), .RSTB(sys_rst_l), .Q(rec_dataH_temp_0_) );
 SDFFARX1 rec_dataH_reg_0_ ( .D(rec_dataH_temp_0_), .SI(xmit_doneH), .SE(test_se), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(rec_dataH[0]) );
 u_xmit_test_1 iXMIT ( .sys_clk(sys_clk), .sys_rst_l(sys_rst_l), .uart_xmitH(uart_XMIT_dataH), .xmitH(xmitH), .xmit_dataH(xmit_dataH), .xmit_doneH(xmit_doneH), .uart_test_mode_in(test_mode), .test_si(n18), .test_se(test_se) );
 u_rec_test_1 iRECEIVER ( .sys_rst_l(sys_rst_l),